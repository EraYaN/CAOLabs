library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity memory is
	port
	(
		clk			: in  std_logic;
		rst			: in  std_logic;
		memread			: in  std_logic;
		memwrite		: in  std_logic;
		address1		: in  std_logic_vector (31 downto 0);
		address2		: in  std_logic_vector (31 downto 0);
		writedata		: in  std_logic_vector (31 downto 0);
		instruction		: out std_logic_vector (31 downto 0);
		readdata		: out std_logic_vector (31 downto 0)
	);
end memory;

architecture behavior of memory is
	type ramcell is array (0 to 255) of std_logic_vector (7 downto 0);
	signal ram			: ramcell;
	signal masked1, masked2		: std_logic_vector (7 downto 0);
	signal selector1, selector2	: natural range 0 to 255;
begin
	masked1 <= address1 (7 downto 2) & "00";
	masked2 <= address2 (7 downto 2) & "00";
	selector1 <= to_integer (unsigned (masked1));
	selector2 <= to_integer (unsigned (masked2));

	process (clk, rst, memread, memwrite, address1, address2, writedata)
	begin
		if (rising_edge (clk)) then
			if (rst = '1') then
				ram (  0) <= "00100101"; -- move $s4,$zero
				ram (  1) <= "10100000";
				ram (  2) <= "00000000";
				ram (  3) <= "00000000";
				ram (  4) <= "00100101"; -- move $s5,$zero
				ram (  5) <= "10101000";
				ram (  6) <= "00000000";
				ram (  7) <= "00000000";
				ram (  8) <= "00010010"; -- addi $t1,$zero,18
				ram (  9) <= "00000000";
				ram ( 10) <= "00001001";
				ram ( 11) <= "00100000";
				ram ( 12) <= "00000100"; -- addi $s0,$zero,4
				ram ( 13) <= "00000000";
				ram ( 14) <= "00010000";
				ram ( 15) <= "00100000";
				ram ( 16) <= "00000001"; -- addi $s2,$zero,1
				ram ( 17) <= "00000000";
				ram ( 18) <= "00010010";
				ram ( 19) <= "00100000";
				ram ( 20) <= "10000000"; -- sll  $s2,$s2,22
				ram ( 21) <= "10010101";
				ram ( 22) <= "00010010";
				ram ( 23) <= "00000000";
				ram ( 24) <= "00101100"; -- addi $s2,$s2,44
				ram ( 25) <= "00000000";
				ram ( 26) <= "01010010";
				ram ( 27) <= "00100010";
				ram ( 28) <= "11111110"; -- addi $s6,$zero,-2
				ram ( 29) <= "11111111";
				ram ( 30) <= "00010110";
				ram ( 31) <= "00100000";
				ram ( 32) <= "00000100"; -- sllv $s0,$s0,$s6
				ram ( 33) <= "10000000";
				ram ( 34) <= "11010000";
				ram ( 35) <= "00000010";
				ram ( 36) <= "00001001"; -- jalr $s1,$s2
				ram ( 37) <= "10001000";
				ram ( 38) <= "01000000";
				ram ( 39) <= "00000010";
				ram ( 40) <= "00001000"; -- addi $s4,$s4,8
				ram ( 41) <= "00000000";
				ram ( 42) <= "10010100";
				ram ( 43) <= "00100010";
				ram ( 44) <= "00001001"; -- addi $s5,$s5,9
				ram ( 45) <= "00000000";
				ram ( 46) <= "10110101";
				ram ( 47) <= "00100010";
				ram ( 48) <= "00000001"; -- beq $s5,$t1,done
				ram ( 49) <= "00000000";
				ram ( 50) <= "10101001";
				ram ( 51) <= "00010010";
				ram ( 52) <= "00001000"; -- jr $s1
				ram ( 53) <= "00000000";
				ram ( 54) <= "00100000";
				ram ( 55) <= "00000010";
				ram ( 56) <= "00000100"; -- done:  sllv $s4,$s4,$s4
				ram ( 57) <= "10100000";
				ram ( 58) <= "10010100";
				ram ( 59) <= "00000010";
				for i in 60 to 255 loop
					ram (i) <= std_logic_vector (to_unsigned (0, 8));
				end loop;
			else
				if (memwrite = '1') then
					ram (selector2 + 0) <= writedata (7 downto 0);
					ram (selector2 + 1) <= writedata (15 downto 8);
					ram (selector2 + 2) <= writedata (23 downto 16);
					ram (selector2 + 3) <= writedata (31 downto 24);
				end if;
			end if;
		end if;
	end process;
	instruction <= ram (selector1 + 3) & ram (selector1 + 2) & ram (selector1 + 1) & ram (selector1 + 0);
	with memread select
		readdata <=	std_logic_vector (to_unsigned (0, 32)) when '0',
				ram (selector2 + 3) & ram (selector2 + 2) & ram (selector2 + 1) & ram (selector2 + 0) when others;
end behavior;
